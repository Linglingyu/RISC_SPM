library verilog;
use verilog.vl_types.all;
entity Control_Unit is
    generic(
        word_size       : integer := 8;
        op_size         : integer := 4;
        state_size      : integer := 4;
        src_size        : integer := 2;
        dest_size       : integer := 2;
        Sel1_size       : integer := 3;
        Sel2_size       : integer := 2;
        S_idle          : integer := 0;
        S_fet1          : integer := 1;
        S_fet2          : integer := 2;
        S_dec           : integer := 3;
        S_ex1           : integer := 4;
        S_rd1           : integer := 5;
        S_rd2           : integer := 6;
        S_wr1           : integer := 7;
        S_wr2           : integer := 8;
        S_br1           : integer := 9;
        S_br2           : integer := 10;
        S_halt          : integer := 11;
        NOP             : integer := 0;
        ADD             : integer := 1;
        SUB             : integer := 2;
        \AND\           : integer := 3;
        \NOT\           : integer := 4;
        RD              : integer := 5;
        WR              : integer := 6;
        BR              : integer := 7;
        BRZ             : integer := 8;
        R0              : integer := 0;
        R1              : integer := 1;
        R2              : integer := 2;
        R3              : integer := 3
    );
    port(
        Load_R0         : out    vl_logic;
        Load_R1         : out    vl_logic;
        Load_R2         : out    vl_logic;
        Load_R3         : out    vl_logic;
        Load_PC         : out    vl_logic;
        Inc_PC          : out    vl_logic;
        Sel_Bus_1_Mux   : out    vl_logic_vector;
        Sel_Bus_2_Mux   : out    vl_logic_vector;
        Load_IR         : out    vl_logic;
        Load_Add_R      : out    vl_logic;
        Load_Reg_Y      : out    vl_logic;
        Load_Reg_Z      : out    vl_logic;
        write           : out    vl_logic;
        instruction     : in     vl_logic_vector;
        zero            : in     vl_logic;
        clk             : in     vl_logic;
        rst             : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of word_size : constant is 1;
    attribute mti_svvh_generic_type of op_size : constant is 1;
    attribute mti_svvh_generic_type of state_size : constant is 1;
    attribute mti_svvh_generic_type of src_size : constant is 1;
    attribute mti_svvh_generic_type of dest_size : constant is 1;
    attribute mti_svvh_generic_type of Sel1_size : constant is 1;
    attribute mti_svvh_generic_type of Sel2_size : constant is 1;
    attribute mti_svvh_generic_type of S_idle : constant is 1;
    attribute mti_svvh_generic_type of S_fet1 : constant is 1;
    attribute mti_svvh_generic_type of S_fet2 : constant is 1;
    attribute mti_svvh_generic_type of S_dec : constant is 1;
    attribute mti_svvh_generic_type of S_ex1 : constant is 1;
    attribute mti_svvh_generic_type of S_rd1 : constant is 1;
    attribute mti_svvh_generic_type of S_rd2 : constant is 1;
    attribute mti_svvh_generic_type of S_wr1 : constant is 1;
    attribute mti_svvh_generic_type of S_wr2 : constant is 1;
    attribute mti_svvh_generic_type of S_br1 : constant is 1;
    attribute mti_svvh_generic_type of S_br2 : constant is 1;
    attribute mti_svvh_generic_type of S_halt : constant is 1;
    attribute mti_svvh_generic_type of NOP : constant is 1;
    attribute mti_svvh_generic_type of ADD : constant is 1;
    attribute mti_svvh_generic_type of SUB : constant is 1;
    attribute mti_svvh_generic_type of \AND\ : constant is 1;
    attribute mti_svvh_generic_type of \NOT\ : constant is 1;
    attribute mti_svvh_generic_type of RD : constant is 1;
    attribute mti_svvh_generic_type of WR : constant is 1;
    attribute mti_svvh_generic_type of BR : constant is 1;
    attribute mti_svvh_generic_type of BRZ : constant is 1;
    attribute mti_svvh_generic_type of R0 : constant is 1;
    attribute mti_svvh_generic_type of R1 : constant is 1;
    attribute mti_svvh_generic_type of R2 : constant is 1;
    attribute mti_svvh_generic_type of R3 : constant is 1;
end Control_Unit;
